module batalha_naval (
    
);
    
endmodule